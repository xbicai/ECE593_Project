`define FIFO_WIDTH	8
`define FIFO_ADDR	2
`define FIFO_DEPTH	2**`FIFO_ADDR