`define FIFO_WIDTH	8
`define FIFO_DEPTH	4