`define UVM_REPORT_DISABLE_FILE_LINE    // removes file line section in uvm_info prints for clarity
`define FIFO_WIDTH	8
`define FIFO_ADDR	2
`define FIFO_DEPTH	2**`FIFO_ADDR
`define SEQ_DELAY_L #500
`define SEQ_DELAY_S #100