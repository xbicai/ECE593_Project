package new_proj_pkg;
  `include "transaction.sv"
  `include "generator.sv"
  `include "driver.sv"
  `include "monitor.sv"
  `include "scoreboard.sv"
  `include "env.sv"
  `include "async_fifo_test.sv"
endpackage
