// `include "transaction.sv"

class async_fifo_scoreboard #(parameter SIZE = 32);
	

	//------------------------------------------------------------
	// Standard UVM Constructor
	//------------------------------------------------------------


endclass : async_fifo_scoreboard