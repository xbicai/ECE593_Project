package new_proj_pkg;
  `include "transaction.sv"
  `include "generator.sv"
  `include "driver.sv"
  `include "monitor_wr.sv"
  `include "monitor_rd.sv"
  `include "scoreboard.sv"
  `include "env.sv"
endpackage
