package class_tb_pkg;
	`include "./class/transaction.sv"
	`include "./class/generator.sv"
	`include "./class/driver.sv"
	`include "./class/monitor.sv"
	`include "./class/scoreboard.sv"
	`include "./class/env.sv"
	`include "./class/test.sv"
endpackage
