`define W_CYCLE   10        // write clock cycle
`define R_CYCLE   15        // read clock cycle
`define CLK_SHIFT 0     
`define DATA 	  8         // DATA of data
`define ADDR 	  4         // amount of addresses
`define DEPTH     2**`ADDR  // how many total addresses