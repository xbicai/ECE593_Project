// `include "env.sv"

class test;

	//------------------------------------------------------------
	// Standard UVM Constructor
	//------------------------------------------------------------


endclass